LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY POS_CONV IS
	PORT(
			LPOS : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			SIZE : IN STD_LOGIC;
			XPOS : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
			YPOS : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
		);
END POS_CONV;

ARCHITECTURE main OF POS_CONV IS
BEGIN
	PROCESS(LPOS, SIZE)
	VARIABLE LP : STD_LOGIC_VECTOR(10 DOWNTO 0);
	VARIABLE SZ : INTEGER RANGE 0 TO 40;
	BEGIN
		IF(SIZE = '0') THEN
			SZ := 40;
		ELSE
			SZ := 20;
		END IF;
		LP := LPOS(10 DOWNTO 0);
		XPOS <= conv_std_logic_vector(conv_integer(LP) MOD SZ, 6);
		YPOS <= conv_std_logic_vector(conv_integer(LP) / SZ, 5);
	END PROCESS;
END main;