LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY ALU IS
	PORT(
			X : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			OP : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			FR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			RES : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
END ALU;

ARCHITECTURE main OF ALU IS
BEGIN
END main;